----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:41:04 01/25/2019 
-- Design Name: 
-- Module Name:    Practicando_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Practicando_1 is
port(S0,S1,S2,S3,S4,S5,S6 : out std_logic;

end Practicando_1;

architecture Behavioral of Practicando_1 is

begin
--Esto es un comentario
S0:=5#123
S1:='A'
S2:=B"0111010001010100001010111010100010101011101010010010100"
S3:=5.15

end Behavioral;

